module ppu();

endmodule